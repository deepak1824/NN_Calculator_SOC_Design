//
// This is a simple interface for the design reset;
//

interface tbRESET(output reg RESET);



endinterface : tbRESET
